//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
`timescale 1ns/1ns
module
UART_UART_0_COREUART
(
RESET_N
,
CLK
,
WEN
,
OEN
,
CSN
,
DATA_IN
,
RX
,
BAUD_VAL
,
BIT8
,
PARITY_EN
,
ODD_N_EVEN
,
PARITY_ERR
,
OVERFLOW
,
TXRDY
,
RXRDY
,
DATA_OUT
,
TX
,
FRAMING_ERR
)
;
parameter
TX_FIFO
=
0
;
parameter
RX_FIFO
=
0
;
parameter
RX_LEGACY_MODE
=
0
;
parameter
FAMILY
=
15
;
input
RESET_N
;
input
CLK
;
input
WEN
;
input
OEN
;
input
CSN
;
input
[
7
:
0
]
DATA_IN
;
input
RX
;
input
[
12
:
0
]
BAUD_VAL
;
input
BIT8
;
input
PARITY_EN
;
input
ODD_N_EVEN
;
output
PARITY_ERR
;
output
OVERFLOW
;
output
TXRDY
;
output
RXRDY
;
output
[
7
:
0
]
DATA_OUT
;
output
TX
;
output
FRAMING_ERR
;
`define S0  \
2 \
'b \
00
`define S1  \
2 \
'b \
01
`define CUARTOOI  \
2 \
'b \
10
`define CUARTIOI  \
2 \
'b \
11
wire
PARITY_ERR
;
wire
FRAMING_ERR
;
wire
OVERFLOW
;
wire
CUARTlOI
;
wire
TXRDY
;
reg
RXRDY
;
wire
CUARTOII
;
wire
CUARTIII
;
wire
CUARTlII
;
reg
[
7
:
0
]
DATA_OUT
;
wire
TX
;
wire
CUARTll
;
wire
CUARTIl
;
wire
CUARTOlI
;
reg
[
7
:
0
]
CUARTIlI
;
wire
[
7
:
0
]
CUARTllI
;
wire
[
7
:
0
]
CUARTO0I
;
wire
CUARTI0I
;
reg
[
7
:
0
]
CUARTl0I
;
wire
[
7
:
0
]
CUARTO1I
;
wire
[
7
:
0
]
CUARTI1I
;
wire
CUARTl1I
;
wire
CUARTOOl
;
reg
CUARTIOl
;
reg
CUARTlOl
;
wire
CUARTOIl
;
wire
CUARTIIl
;
wire
CUARTlIl
;
wire
CUARTOll
;
wire
CUARTIll
;
wire
CUARTlll
;
reg
CUARTO0l
;
reg
CUARTI0l
;
wire
CUARTl0l
;
reg
CUARTO1l
;
reg
CUARTI1l
;
reg
CUARTl1l
;
reg
CUARTOO0
;
reg
CUARTIO0
;
reg
CUARTlO0
;
reg
[
1
:
0
]
CUARTOI0
;
reg
[
1
:
0
]
CUARTII0
;
wire
CUARTlI0
;
wire
CUARTOl0
;
reg
CUARTIl0
;
wire
CUARTll0
;
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
:
CUARTO00
if
(
RESET_N
==
1
'b
0
)
begin
CUARTIlI
<=
{
8
{
1
'b
0
}
}
;
CUARTlOl
<=
1
'b
1
;
end
else
begin
CUARTlOl
<=
1
'b
1
;
if
(
CSN
==
1
'b
0
&
WEN
==
1
'b
0
)
begin
CUARTIlI
<=
DATA_IN
;
CUARTlOl
<=
1
'b
0
;
end
end
end
assign
CUARTOlI
=
WEN
==
1
'b
0
&
CSN
==
1
'b
0
?
1
'b
1
:
1
'b
0
;
always
@
(
CUARTO1I
or
CUARTl0I
or
PARITY_ERR
)
begin
if
(
RX_FIFO
==
1
'b
0
)
begin
DATA_OUT
=
CUARTO1I
;
end
else
begin
if
(
PARITY_ERR
==
1
'b
1
)
begin
DATA_OUT
=
CUARTO1I
;
end
else
begin
DATA_OUT
=
CUARTl0I
;
end
end
end
assign
CUARTI0I
=
(
RX_FIFO
==
1
'b
0
)
?
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
)
:
!
CUARTlIl
;
assign
CUARTOll
=
(
RX_FIFO
==
1
'b
0
)
?
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
)
:
CUARTI0l
;
assign
CUARTIll
=
(
RX_FIFO
==
1
'b
0
)
?
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
)
:
CUARTI1l
;
assign
CUARTll0
=
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
;
assign
CUARTI1I
=
(
PARITY_ERR
==
1
'b
0
)
?
CUARTO1I
:
8
'b
0
;
generate
if
(
RX_LEGACY_MODE
==
1
'b
1
)
begin
always
@
(
CUARTOII
or
CUARTIO0
)
begin
if
(
RX_FIFO
==
1
'b
0
)
begin
RXRDY
=
CUARTOII
;
end
else
begin
RXRDY
=
!
CUARTIO0
;
end
end
end
else
begin
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
RXRDY
=
1
'b
0
;
end
else
begin
if
(
RX_FIFO
==
1
'b
0
)
begin
if
(
CUARTlI0
==
1
'b
1
||
CUARTOII
==
1
'b
0
)
begin
RXRDY
=
CUARTOII
;
end
end
else
begin
if
(
CUARTlI0
==
1
'b
1
||
(
CUARTIO0
==
1
'b
1
)
||
(
(
CUARTIO0
==
1
'b
0
)
&&
(
CUARTOl0
==
1
'b
1
)
)
)
begin
RXRDY
=
!
CUARTIO0
;
end
end
end
end
end
endgenerate
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
CUARTI0l
<=
1
'b
0
;
CUARTO0l
<=
1
'b
0
;
end
else
begin
CUARTO0l
<=
CUARTlll
;
CUARTI0l
<=
CUARTO0l
;
end
end
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
CUARTI1l
<=
1
'b
0
;
CUARTO1l
<=
1
'b
0
;
end
else
begin
CUARTO1l
<=
CUARTl0l
;
CUARTI1l
<=
CUARTO1l
;
end
end
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
CUARTOI0
<=
`S0
;
end
else
begin
CUARTOI0
<=
CUARTII0
;
end
end
always
@
(
CUARTOI0
,
CUARTIO0
,
CUARTOOl
)
begin
CUARTII0
=
CUARTOI0
;
CUARTIOl
=
1
'b
1
;
CUARTl1l
=
1
'b
0
;
case
(
CUARTOI0
)
`S0
:
if
(
CUARTIO0
==
1
'b
1
&&
CUARTOOl
==
1
'b
0
)
begin
CUARTII0
=
`S1
;
CUARTIOl
=
1
'b
0
;
end
`S1
:
CUARTII0
=
`CUARTOOI
;
`CUARTOOI
:
CUARTII0
=
`CUARTIOI
;
`CUARTIOI
:
begin
CUARTII0
=
`S0
;
CUARTl1l
=
1
'b
1
;
end
endcase
end
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
CUARTl0I
<=
{
8
{
1
'b
0
}
}
;
end
else
begin
if
(
CUARTl1l
==
1
'b
1
)
begin
CUARTl0I
<=
CUARTO0I
;
end
end
end
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
CUARTIO0
<=
1
'b
1
;
CUARTlO0
<=
1
'b
1
;
end
else
begin
if
(
CUARTl1l
==
1
'b
1
)
begin
CUARTIO0
<=
1
'b
0
;
end
else
begin
if
(
CSN
==
1
'b
0
&&
OEN
==
1
'b
0
)
begin
CUARTIO0
<=
1
'b
1
;
end
end
CUARTlO0
<=
CUARTIO0
;
end
end
always
@
(
posedge
CLK
or
negedge
RESET_N
)
begin
if
(
RESET_N
==
1
'b
0
)
begin
CUARTIl0
<=
1
'b
0
;
end
else
begin
if
(
CUARTlII
==
1
'b
0
&&
CUARTlIl
==
1
'b
1
)
CUARTIl0
<=
1
'b
1
;
else
if
(
CUARTll0
==
1
'b
1
)
CUARTIl0
<=
1
'b
0
;
else
CUARTIl0
<=
CUARTIl0
;
end
end
assign
OVERFLOW
=
(
RX_FIFO
==
1
'b
0
)
?
CUARTlOI
:
CUARTIl0
;
assign
CUARTIII
=
(
(
PARITY_ERR
==
1
'b
1
)
||
CUARTlIl
==
1
'b
1
)
?
1
'b
1
:
CUARTlII
;
UART_UART_0_Clock_gen
CUARTI00
(
.CUARTII
(
CLK
)
,
.CUARTlI
(
RESET_N
)
,
.CUARTOl
(
BAUD_VAL
)
,
.CUARTIl
(
CUARTIl
)
,
.CUARTll
(
CUARTll
)
)
;
UART_UART_0_Tx_async
#
(
.TX_FIFO
(
TX_FIFO
)
)
CUARTl00
(
.CUARTII
(
CLK
)
,
.CUARTll
(
CUARTll
)
,
.CUARTlI
(
RESET_N
)
,
.CUARTOlI
(
CUARTOlI
)
,
.CUARTIlI
(
CUARTIlI
)
,
.CUARTllI
(
CUARTllI
)
,
.CUARTO10
(
CUARTl1I
)
,
.CUARTI10
(
CUARTIIl
)
,
.CUARTl10
(
BIT8
)
,
.CUARTOO1
(
PARITY_EN
)
,
.CUARTIO1
(
ODD_N_EVEN
)
,
.CUARTlO1
(
TXRDY
)
,
.CUARTOI1
(
TX
)
,
.CUARTOIl
(
CUARTOIl
)
)
;
UART_UART_0_Rx_async
#
(
.RX_FIFO
(
RX_FIFO
)
,
.RX_LEGACY_MODE
(
RX_LEGACY_MODE
)
)
CUARTII1
(
.CUARTII
(
CLK
)
,
.CUARTIl
(
CUARTIl
)
,
.CUARTlI
(
RESET_N
)
,
.CUARTl10
(
BIT8
)
,
.CUARTOO1
(
PARITY_EN
)
,
.CUARTIO1
(
ODD_N_EVEN
)
,
.CUARTI0I
(
CUARTI0I
)
,
.CUARTOll
(
CUARTOll
)
,
.CUARTlI1
(
FRAMING_ERR
)
,
.CUARTIll
(
CUARTIll
)
,
.CUARTlI0
(
CUARTlI0
)
,
.CUARTOl0
(
CUARTOl0
)
,
.CUARTOl1
(
RX
)
,
.CUARTIl1
(
CUARTlOI
)
,
.CUARTll1
(
PARITY_ERR
)
,
.CUARTlll
(
CUARTlll
)
,
.CUARTl0l
(
CUARTl0l
)
,
.CUARTOII
(
CUARTOII
)
,
.CUARTO1I
(
CUARTO1I
)
,
.CUARTlII
(
CUARTlII
)
)
;
generate
if
(
TX_FIFO
==
1
'b
1
)
begin
UART_UART_0_fifo_256x8
CUARTO01
(
.CUARTI01
(
CUARTllI
)
,
.CUARTl01
(
CLK
)
,
.CUARTO11
(
CLK
)
,
.CUARTI11
(
CUARTIlI
)
,
.WRB
(
CUARTlOl
)
,
.RDB
(
CUARTOIl
)
,
.RESET
(
RESET_N
)
,
.FULL
(
CUARTIIl
)
,
.EMPTY
(
CUARTl1I
)
)
;
end
endgenerate
generate
if
(
RX_FIFO
==
1
'b
1
)
begin
UART_UART_0_fifo_256x8
CUARTl11
(
.CUARTI01
(
CUARTO0I
)
,
.CUARTl01
(
CLK
)
,
.CUARTO11
(
CLK
)
,
.CUARTI11
(
CUARTI1I
)
,
.WRB
(
CUARTIII
)
,
.RDB
(
CUARTIOl
)
,
.RESET
(
RESET_N
)
,
.FULL
(
CUARTlIl
)
,
.EMPTY
(
CUARTOOl
)
)
;
end
endgenerate
endmodule
