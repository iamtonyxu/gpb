`timescale 1ns/100ps

module CORECAN_wrapper
(
    // OPB Interface
    input               OPB_CLK,
    input               OPB_RST,
    input      [10:0]   OPB_ADDR,
    input      [31:0]   OPB_DI,
    output     [31:0]   OPB_DO,
    input               OPB_WE,
    input               OPB_RE,

    // CAN Interface
    output              CAN_TX_EN_N,
    output              CAN_TX,
    input               CAN_RX

);

// apb bus signals
wire pclk, presetn, psel;
wire pwrite; // OPB_WE driven, and it will last two cycles
wire penable; // It goes after OPB_RE or OPB_WE, and will last one cycle
reg [10:0] paddr; // 11 bits address, from OPB_ADDR[10:0]
reg [31:0] pwdata; // from OPB_DI[31:0]
wire [31:0] prdata; // to OPB_DO[31:0]

// OPB to APB signal conversion
assign pclk = OPB_CLK; // 100MHz clock
assign presetn = ~OPB_RST;
assign psel = 1'b1; // always selected
assign OPB_DO = prdata; // APB read data to OPB read data

// latch address and write data at OPB_CLK rising edge
always @(posedge OPB_CLK or posedge OPB_RST) begin
    if (OPB_RST) begin
        paddr <= 11'b0;
        pwdata <= 32'b0;
    end else if (OPB_WE || OPB_RE) begin
        paddr <= OPB_ADDR[10:0];
        pwdata <= OPB_DI[31:0];
    end
end

// pwrite lasts two cycles, penable lasts one cycle
reg pwrite_d1, pwrite_d2;
always @(posedge OPB_CLK or posedge OPB_RST) begin
    if (OPB_RST) begin
        pwrite_d1 <= 1'b0;
        pwrite_d2 <= 1'b0;
    end else begin
        pwrite_d1 <= OPB_WE;
        pwrite_d2 <= pwrite_d1;
    end
end

// pread lasts two cycles, penable lasts one cycle
reg pread_d1, pread_d2;
always @(posedge OPB_CLK or posedge OPB_RST) begin
    if (OPB_RST) begin
        pread_d1 <= 1'b0;
        pread_d2 <= 1'b0;
    end else begin
        pread_d1 <= OPB_RE;
        pread_d2 <= pread_d1;
    end
end

assign pwrite = pwrite_d1 || pwrite_d2;
assign penable = pwrite_d2 || pread_d2;

// Instantiate the CORECAN module
CORECAN_C0 uut (
    // APB Interface
    .PCLK(pclk),
    .PRESETN(presetn),
    .PSEL(psel),
    .PENABLE(penable),
    .PWRITE(pwrite),
    .PADDR(paddr),
    .PWDATA(pwdata),
    .PRDATA(prdata),
    .PREADY(), // Always ready in this example
    .INT_N(), // Interrupt not used in this example

    // CAN Interface
    .CAN_TX_EN_N(CAN_TX_EN_N),
    .CAN_TX(CAN_TX),
    .CAN_RX(CAN_RX)
);

endmodule


/*
// CoreCan IP generated by Libero
module CORECAN_C0(
    // APB Interface
    input PCLK,
    input PRESETN,
    input PSEL,
    input PENABLE,
    input PWRITE,
    input [10:0] PADDR,
    input [31:0] PWDATA,
    output [31:0] PRDATA,
    output PREADY,
    output INT_N,

    // CAN Interface
    output CAN_TX_EN_N,
    output CAN_TX,
    input CAN_RX
);
*/