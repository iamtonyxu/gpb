//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
`timescale 1ns/1ns
module
UART_UART_0_Tx_async
(
CUARTII
,
CUARTll
,
CUARTlI
,
CUARTOlI
,
CUARTIlI
,
CUARTllI
,
CUARTO10
,
CUARTI10
,
CUARTl10
,
CUARTOO1
,
CUARTIO1
,
CUARTlO1
,
CUARTOI1
,
CUARTOIl
)
;
parameter
TX_FIFO
=
0
;
input
CUARTII
;
input
CUARTll
;
input
CUARTlI
;
input
CUARTOlI
;
input
[
7
:
0
]
CUARTIlI
;
input
[
7
:
0
]
CUARTllI
;
input
CUARTO10
;
input
CUARTI10
;
input
CUARTl10
;
input
CUARTOO1
;
input
CUARTIO1
;
output
CUARTlO1
;
wire
CUARTlO1
;
output
CUARTOI1
;
output
CUARTOIl
;
reg
CUARTOI1
;
parameter
CUARTllIl
=
0
;
parameter
CUARTO0Il
=
1
;
parameter
CUARTI0Il
=
2
;
parameter
CUARTl0Il
=
3
;
parameter
CUARTO1Il
=
4
;
parameter
CUARTI1Il
=
5
;
parameter
CUARTl1Il
=
6
;
integer
CUARTOOll
;
reg
CUARTIOll
;
reg
[
7
:
0
]
CUARTlOll
;
reg
[
3
:
0
]
CUARTOIll
;
reg
CUARTIIll
;
wire
CUARTOIl
;
reg
CUARTlIll
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOlll
if
(
!
CUARTlI
)
begin
CUARTIOll
<=
1
'b
1
;
end
else
begin
if
(
TX_FIFO
==
1
'b
0
)
begin
if
(
CUARTll
)
begin
if
(
CUARTOOll
==
CUARTI0Il
)
begin
CUARTIOll
<=
1
'b
1
;
end
end
if
(
CUARTOlI
)
begin
CUARTIOll
<=
1
'b
0
;
end
end
else
begin
CUARTIOll
<=
!
CUARTI10
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTIlll
if
(
!
CUARTlI
)
begin
CUARTOOll
<=
CUARTllIl
;
CUARTlOll
<=
8
'b
0
;
CUARTlIll
<=
1
'b
1
;
end
else
begin
if
(
CUARTll
||
(
CUARTOOll
==
CUARTllIl
)
||
(
CUARTOOll
==
CUARTl1Il
)
||
(
CUARTOOll
==
CUARTO0Il
)
)
begin
CUARTlIll
<=
1
'b
1
;
case
(
CUARTOOll
)
CUARTllIl
:
begin
if
(
TX_FIFO
==
1
'b
0
)
begin
if
(
!
CUARTIOll
)
begin
CUARTOOll
<=
CUARTO0Il
;
end
else
begin
CUARTOOll
<=
CUARTllIl
;
end
end
else
begin
if
(
CUARTO10
==
1
'b
0
)
begin
CUARTlIll
<=
1
'b
0
;
CUARTOOll
<=
CUARTl1Il
;
end
else
begin
CUARTOOll
<=
CUARTllIl
;
CUARTlIll
<=
1
'b
1
;
end
end
end
CUARTO0Il
:
begin
CUARTOOll
<=
CUARTI0Il
;
end
CUARTI0Il
:
begin
CUARTOOll
<=
CUARTl0Il
;
if
(
TX_FIFO
==
1
'b
0
)
begin
CUARTlOll
<=
CUARTIlI
;
end
else
begin
CUARTlOll
<=
CUARTllI
;
end
end
CUARTl0Il
:
begin
if
(
CUARTl10
)
begin
if
(
CUARTOIll
==
4
'b
0111
)
begin
if
(
CUARTOO1
)
begin
CUARTOOll
<=
CUARTO1Il
;
end
else
begin
CUARTOOll
<=
CUARTI1Il
;
end
end
else
begin
CUARTOOll
<=
CUARTl0Il
;
end
end
else
begin
if
(
CUARTOIll
==
4
'b
0110
)
begin
if
(
CUARTOO1
)
begin
CUARTOOll
<=
CUARTO1Il
;
end
else
begin
CUARTOOll
<=
CUARTI1Il
;
end
end
else
begin
CUARTOOll
<=
CUARTl0Il
;
end
end
end
CUARTO1Il
:
begin
CUARTOOll
<=
CUARTI1Il
;
end
CUARTI1Il
:
begin
CUARTOOll
<=
CUARTllIl
;
end
CUARTl1Il
:
begin
CUARTOOll
<=
CUARTO0Il
;
end
default
:
begin
CUARTOOll
<=
CUARTllIl
;
end
endcase
end
end
end
assign
CUARTOIl
=
CUARTlIll
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTllll
if
(
!
CUARTlI
)
begin
CUARTOIll
<=
4
'b
0000
;
end
else
begin
if
(
CUARTll
)
begin
if
(
CUARTOOll
!=
CUARTl0Il
)
begin
CUARTOIll
<=
4
'b
0000
;
end
else
begin
CUARTOIll
<=
CUARTOIll
+
1
'b
1
;
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTO0ll
if
(
!
CUARTlI
)
begin
CUARTOI1
<=
1
'b
1
;
end
else
begin
if
(
CUARTll
||
(
CUARTOOll
==
CUARTllIl
)
||
(
CUARTOOll
==
CUARTl1Il
)
||
(
CUARTOOll
==
CUARTO0Il
)
)
begin
case
(
CUARTOOll
)
CUARTllIl
:
begin
CUARTOI1
<=
1
'b
1
;
end
CUARTO0Il
:
begin
CUARTOI1
<=
1
'b
1
;
end
CUARTI0Il
:
begin
CUARTOI1
<=
1
'b
0
;
end
CUARTl0Il
:
begin
CUARTOI1
<=
CUARTlOll
[
CUARTOIll
]
;
end
CUARTO1Il
:
begin
CUARTOI1
<=
CUARTIO1
^
CUARTIIll
;
end
CUARTI1Il
:
begin
CUARTOI1
<=
1
'b
1
;
end
default
:
begin
CUARTOI1
<=
1
'b
1
;
end
endcase
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTI0ll
if
(
!
CUARTlI
)
begin
CUARTIIll
<=
1
'b
0
;
end
else
begin
if
(
CUARTll
&
CUARTOO1
)
begin
if
(
CUARTOOll
==
CUARTl0Il
)
begin
CUARTIIll
<=
CUARTIIll
^
CUARTlOll
[
CUARTOIll
]
;
end
else
begin
CUARTIIll
<=
CUARTIIll
;
end
end
if
(
CUARTOOll
==
CUARTI1Il
)
begin
CUARTIIll
<=
1
'b
0
;
end
end
end
assign
CUARTlO1
=
CUARTIOll
;
endmodule
