`timescale 1ns/100ps
/*
* File: cmn_pwm_wrapper.v
*
* Description:
*
*   This module is a wrapper for the cmn_pwm module. It connects the OPB interface to the cmn_pwm module.
*   It also includes the necessary clock and reset signals.
*   1. OPB Write mot_pwm_param01/23/45 or brk_pwm_param
*   2. OPB Read mot_pwm_param01/23/45 or brk_pwm_param and check
*   3. OPB Write pwm_config to select test mode and enable/disable PWM
*   4. OPB Read pwm_config to check test mode and enable/disable PWM
*   5. OPB Write pwm_start to start PWM generation
*   6. OPB Read pwm_status if need
*
*/

`define ADDR_PWM_CONFIG         4'h0
`define ADDR_MOT_PWM_PARAM01    4'h1
`define ADDR_MOT_PWM_PARAM23    4'h2
`define ADDR_MOT_PWM_PARAM45    4'h3
`define ADDR_BRK_PWM_PARAM      4'h4
`define ADDR_PWM_CONTROL        4'h5
`define ADDR_PWM_STATUS         4'h6

module cmn_pwm_wrapper
(
    // OPB signals
    input                   OPB_CLK,        // 100MHz clock
    input                   OPB_RST,        // Reset signal
    input                   OPB_RE,         // OPB read enable
    input                   OPB_WE,         // OPB write enable
    input       [31:0]      OPB_ADDR,       // OPB address bus
    output reg  [31:0]      OPB_DO,         // OPB data output
    input       [31:0]      OPB_DI,         // OPB data input

    // Motor and brake signals
    output      [5:0]       mot_pwm_o,      // Motor PWM output
    output      [1:0]       brk_pwm_o,      // Brake PWM output
    output                  mot_en_out_o,   // Motor enable output
    output                  brk_en_out_o,   // Brake enable output
    input                   mot_over_curr_i,// Motor over-current input
    input                   brk_over_curr_i, // Brake over-current input
    output                  pwm_override_o // 1: override, 0: normal operation
);

    parameter MAX_CNTR_200US = 5000; // 200us at 25MHz
    parameter DEFAULT_TEST_DURATION = 16'd4000; // 100ms at start_pwm_period_out (25us) if test_mode = 1
    parameter MAX_TEST_DURATION = 16'd5000; // 125ms at start_pwm_period_out (25us) if test_mode = 1
    parameter MAX_SYNC_CNTR = 3; // 3 clock cycles at 25MHz
    parameter DEBOUNCE_TIME = 8; // 8 clock cycles  at 25MHz

    // Internal registers
    // pwm_config[2] -> test_mode
    // pwm_config[1] -> mot_pwm_enable
    // pwm_config[0] -> brk_pwm_enable
    // pwm_config[23:8] -> set_test_duration
    reg [31:0] pwm_config;
    // test_mode = 0, free run, FPGA just generate PWM signal without checking over-current signal
    // test_mode = 1, oc-protect mode, FPGA will check over-current signal and stop PWM signal if over-current detected
    wire test_mode; // 0: free-run, 1: oc-protect mode
    wire mot_pwm_enable; // 0: disable, 1: enable
    wire brk_pwm_enable; // 0: disable, 1: enable
    wire [15:0] set_test_duration; // default is 100ms, only used in test_mode = 1

    // mot_pwm_param01, mot_pwm_param23, mot_pwm_param45, brk_pwm_param
    // MOT_PWM_MAX = CLK_RATE_MHZ * 25 * RESOLUTION / 2 - 1 = 25 * 25 * 1 / 2 - 1 = 311
    reg [31:0] mot_pwm_param01; //only [9:0] is used, max value is 311
    reg [31:0] mot_pwm_param23; //only [9:0] is used, max value is 311
    reg [31:0] mot_pwm_param45; //only [9:0] is used, max value is 311
    reg [31:0] brk_pwm_param; //only [9:0] is used, max value is 311
    // pwm_control[0] -> pwm_start, write 1 to start PWM generation and self-clear to 0
    // pwm_control[1] -> pwm_stop, write 1 to stop PWM generation and self-clear to 0
    reg [31:0]pwm_control; // only [1:0] is used
    wire pwm_start; // 0: stop, 1: start
    wire pwm_stop; // 0: stop, 1: stop

    reg [31:0]pwm_status; // pwm_status will be reset if pwm_start = 1
    // pwm_status[0] <- mot_over_curr
    // pwm_status[1] <- brk_over_curr
    // pwm_status[2] <- mot_over_curr_protected
    // pwm_status[3] <- brk_over_curr_protected
    // pwm_status[23:8] <- act_test_duration

    reg [15:0] act_test_duration; // actual test duration, the resolution is 25us, only used in test_mode = 1
    wire start_pwm_period_out; // generated by cmn_pwm, the period is 25us, used to update act_test_duration in test_mode = 1

    // clk_25MHz and pulse_200us
    wire clk_25MHz;
    wire pulse_200us;
    reg [15:0] pulse_200us_cntr;

    // sync signal, 3 clock cycles at 25MHz
    wire sync;
    reg [7:0] sync_cntr;

    // cmn_pwm output signals
    wire [5:0] mot_pwm;
    wire [1:0] brk_pwm;
    wire mot_en_out;
    wire brk_en_out;

    wire filt_mot_over_curr; // filtered motor over-current signal
    wire filt_brk_over_curr; // filtered brake over-current signal

    // OPB write operation
    // pwm_config
    always @(posedge OPB_CLK or posedge OPB_RST) begin
        if (OPB_RST) begin
            pwm_config <= {8'h00, DEFAULT_TEST_DURATION, 8'h00};
        end else if (OPB_WE && OPB_ADDR[3:0] == `ADDR_PWM_CONFIG) begin
            pwm_config <= OPB_DI;
            if(pwm_config[23:8] > MAX_TEST_DURATION) begin
                pwm_config[23:8] <= MAX_TEST_DURATION; // set test duration to max value if it exceeds the limit
            end
        end
    end

    // mot_pwm_param01, mot_pwm_param23, mot_pwm_param45, brk_pwm_param
    always @(posedge OPB_CLK or posedge OPB_RST) begin
        if (OPB_RST) begin
            mot_pwm_param01 <= 0;
            mot_pwm_param23 <= 0;
            mot_pwm_param45 <= 0;
            brk_pwm_param <= 0;
        end else if (OPB_WE && OPB_ADDR[3:0] == `ADDR_MOT_PWM_PARAM01) begin
            mot_pwm_param01 <= OPB_DI;
        end else if (OPB_WE && OPB_ADDR[3:0] == `ADDR_MOT_PWM_PARAM23) begin
            mot_pwm_param23 <= OPB_DI;
        end else if (OPB_WE && OPB_ADDR[3:0] == `ADDR_MOT_PWM_PARAM45) begin
            mot_pwm_param45 <= OPB_DI;
        end else if (OPB_WE && OPB_ADDR[3:0] == `ADDR_BRK_PWM_PARAM) begin
            brk_pwm_param <= OPB_DI;
        end else begin
            mot_pwm_param01 <= mot_pwm_param01;
            mot_pwm_param23 <= mot_pwm_param23;
            mot_pwm_param45 <= mot_pwm_param45;
            brk_pwm_param <= brk_pwm_param;
        end
    end

    // pwm_control
    always @(posedge OPB_CLK or posedge OPB_RST) begin
        if (OPB_RST) begin
            pwm_control <= 0;
        end else if (OPB_WE && OPB_ADDR[3:0] == `ADDR_PWM_CONTROL) begin
            pwm_control <= OPB_DI;
        end else begin
            pwm_control <= 0; // self-clear to 0
        end
    end

    // OPB read operation
    always @(posedge OPB_CLK or posedge OPB_RST) begin
        if (OPB_RST) begin
            OPB_DO <= 0;
        end else if (OPB_RE) begin
            case (OPB_ADDR[3:0])
                `ADDR_PWM_CONFIG: OPB_DO <= pwm_config;
                `ADDR_MOT_PWM_PARAM01: OPB_DO <= mot_pwm_param01;
                `ADDR_MOT_PWM_PARAM23: OPB_DO <= mot_pwm_param23;
                `ADDR_MOT_PWM_PARAM45: OPB_DO <= mot_pwm_param45;
                `ADDR_BRK_PWM_PARAM: OPB_DO <= brk_pwm_param;
                `ADDR_PWM_CONTROL: OPB_DO <= pwm_control;
                `ADDR_PWM_STATUS: OPB_DO <= pwm_status;
                default: OPB_DO <= 0;
            endcase
        end else begin
            OPB_DO <= 0;
        end
    end

    // pwm_config
    assign test_mode = pwm_config[2] ? 1 : 0; // 0: free-run, 1: oc-protect mode
    assign mot_pwm_enable = pwm_config[1] ? 1 : 0; // 0: disable, 1: enable
    assign brk_pwm_enable = pwm_config[0] ? 1 : 0; // 0: disable, 1: enable
    assign set_test_duration = pwm_config[23:8]; // default is 100ms, only used in test_mode = 1

    // pwm_start
    assign pwm_start = pwm_control[0] ? 1 : 0; // 0: stop, 1: start
    // pwm_stop
    assign pwm_stop = pwm_control[1] ? 1 : 0; // 0: stop, 1: stop

    /* state machine
    *
    * ST_IDLE: PWM confguration, and wait for OPB write
    * ST_SYNC: set SYNC singal at least two clock cycles, then go to ST_PWM if pulse_200us = 1
    * ST_PWM: enable PWM output, and align the PWM signal with start_pwm_period_out signal
    * pwm_start will trigger the state from ST_IDLE to ST_PWM when
    * 1) pwm_start = 1 and pwm_stop = 0
    * pwm_start will trigger the state from ST_IDLE to ST_PWM when
    * With test_mode = 0: 
    *   1) pwm_stop = 1; 2) over-current detected
    * With test_mode = 1:
    *   1) pwm_stop = 1;  or 2) after 100ms;  or 3) over-current detected 
    *
    */
    localparam ST_IDLE = 2'b00;
    localparam ST_SYNC = 2'b01;
    localparam ST_PWM = 2'b10;
    reg [1:0] state = ST_IDLE;

    // state machine
    always @(posedge OPB_CLK or posedge OPB_RST) begin
        if (OPB_RST) begin
            state <= ST_IDLE;
        end else begin
            case (state)
                ST_IDLE: begin
                    if (pwm_start) begin
                        state <= ST_SYNC;
                    end else if (pwm_stop) begin
                        state <= ST_IDLE;
                    end else begin
                        state <= ST_IDLE;
                    end
                end
                ST_SYNC: begin
                    if ((sync_cntr >= MAX_SYNC_CNTR) && pulse_200us) begin
                        state <= ST_PWM;
                    end else begin
                        state <= ST_SYNC;
                    end
                end
                ST_PWM: begin
                    if(pwm_stop) begin
                        state <= ST_IDLE;
                    end else if(test_mode) begin
                        if ((act_test_duration == set_test_duration + 1) || filt_mot_over_curr || filt_brk_over_curr) begin
                            state <= ST_IDLE;
                        end else begin
                            state <= ST_PWM;
                        end
                    end else begin
                        if (filt_mot_over_curr || filt_brk_over_curr) begin
                            state <= ST_IDLE; // stop PWM generation if over-current detected
                        end else begin
                            state <= ST_PWM; // continue PWM generation
                        end
                    end
                end
                default: state <= ST_IDLE;
            endcase
        end
    end

    // sync_cntr
    always @(posedge clk_25MHz or posedge OPB_RST) begin
        if (OPB_RST) begin
            sync_cntr <= 0;
        end else if (state == ST_SYNC) begin
            if(sync_cntr < MAX_SYNC_CNTR) begin 
                sync_cntr <= sync_cntr + 1;
            end
        end else if (state == ST_IDLE) begin
            sync_cntr <= 0;
        end
    end

    // act_test_duration
    always @(posedge clk_25MHz or posedge OPB_RST) begin
        if (OPB_RST) begin
            act_test_duration <= 0;
        end else if ((test_mode == 1) && (state == ST_PWM) && start_pwm_period_out) begin
            act_test_duration <= act_test_duration + 1;
        end else if (state == ST_IDLE) begin
            act_test_duration <= 0;
        end
    end

    // pwm_status
    always @(posedge OPB_CLK or posedge OPB_RST) begin
        if (OPB_RST) begin
            pwm_status <= 0;
        end else if(state == ST_PWM) begin
            pwm_status[23:8] <= act_test_duration;
            if(filt_mot_over_curr) begin
                pwm_status[0] <= 1; // over-current detected
            end
            if(filt_brk_over_curr) begin
                pwm_status[1] <= 1; // over-current detected
            end
        end else if (state == ST_IDLE && pwm_start) begin
            pwm_status <= 0; // reset pwm_stat
        end
    end


    // clk_25MHz generation
    CLOCK_DIV clk_16khz_div(
        .CLK_DIV(2),
        .CLK_IN(OPB_CLK),
        .CLK_OUT(clk_25MHz),
        .RST(OPB_RST)
    );

    // pulse_200us generation
    always @(posedge clk_25MHz or posedge OPB_RST) begin
        if (OPB_RST) begin
            pulse_200us_cntr <= 0;
        end else if (pulse_200us_cntr == MAX_CNTR_200US) begin
            pulse_200us_cntr <= 0;
        end else begin
            pulse_200us_cntr <= pulse_200us_cntr + 1;
        end
    end
    assign pulse_200us = (pulse_200us_cntr == MAX_CNTR_200US) ? 1 : 0; // 200us pulse width at 25MHz

     // sync signal, 3 clock cycles at 25MHz
    assign sync = (state == ST_SYNC) && (sync_cntr < MAX_SYNC_CNTR);

    // Instantiate the Unit Under Test (UUT)
    cmn_pwm pwm_0 (
        .reset(OPB_RST),
        .clk(clk_25MHz),
        .sync(sync),
        .pulse_200us(pulse_200us),
        .mot_pwm(mot_pwm),
        .brk_pwm(brk_pwm),
        .mot_en_out(mot_en_out),
        .brk_en_out(brk_en_out),
        .mot_over_curr(mot_over_curr_i),
        .brk_over_curr(brk_over_curr_i),
        .mot_pwm_param01(mot_pwm_param01[9:0]),
        .mot_pwm_param23(mot_pwm_param23[9:0]),
        .mot_pwm_param45(mot_pwm_param45[9:0]),
        .brk_pwm_param(brk_pwm_param[9:0]),
        .mot_en_in(mot_pwm_enable),
        .brk_en_in(brk_pwm_enable),
        .mel_ctrl(1'b1),
        .start_pwm_period_out(start_pwm_period_out)
    );

    // Motor over-current debouncer
    cmn_debouncer #(
        .DEBOUNCE_TIME_LTOH(DEBOUNCE_TIME),
        .DEBOUNCE_TIME_HTOL(DEBOUNCE_TIME)
    ) i_mot_filt (
        .clk(clk_25MHz),
        .reset(OPB_RST),
        .clk_en(1'b1),
        .bypass(1'b0),
        .sig_in(mot_over_curr_i),
        .sig_out(filt_mot_over_curr)
    );

    // Brake over-current debouncer
    cmn_debouncer #(
        .DEBOUNCE_TIME_LTOH(DEBOUNCE_TIME),
        .DEBOUNCE_TIME_HTOL(DEBOUNCE_TIME)
    ) i_brk_filt (
        .clk(clk_25MHz),
        .reset(OPB_RST),
        .clk_en(1'b1),
        .bypass(1'b0),
        .sig_in(brk_over_curr_i),
        .sig_out(filt_brk_over_curr)
    );

    // assign outputs
    assign pwm_override_o = test_mode ? ((state == ST_PWM) && (act_test_duration>0)) : (state == ST_PWM);
    assign mot_pwm_o = (pwm_override_o) ? mot_pwm : 6'b0;
    assign brk_pwm_o = (pwm_override_o) ? brk_pwm : 2'b0;
    assign mot_en_out_o = (pwm_override_o) ? mot_en_out : 1'b0;
    assign brk_en_out_o = (pwm_override_o) ? brk_en_out : 1'b0;

endmodule
