//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
`timescale 1ns/1ns
module
UART_UART_0_Rx_async
(
CUARTII
,
CUARTIl
,
CUARTlI
,
CUARTl10
,
CUARTOO1
,
CUARTIO1
,
CUARTI0I
,
CUARTOll
,
CUARTOl1
,
CUARTIl1
,
CUARTll1
,
CUARTlll
,
CUARTOII
,
CUARTO1I
,
CUARTlII
,
CUARTlI1
,
CUARTIll
,
CUARTl0l
,
CUARTlI0
,
CUARTOl0
)
;
parameter
RX_FIFO
=
0
;
parameter
RX_LEGACY_MODE
=
0
;
input
CUARTII
;
input
CUARTIl
;
input
CUARTlI
;
input
CUARTl10
;
input
CUARTOO1
;
input
CUARTIO1
;
input
CUARTI0I
;
input
CUARTOll
;
input
CUARTIll
;
input
CUARTOl1
;
output
CUARTIl1
;
output
CUARTll1
;
output
CUARTlll
;
output
CUARTOII
;
output
[
7
:
0
]
CUARTO1I
;
output
CUARTlII
;
output
CUARTlI1
;
output
CUARTl0l
;
output
CUARTlI0
;
output
CUARTOl0
;
reg
CUARTlI1
;
reg
CUARTlI0
;
reg
CUARTIl1
;
reg
CUARTll1
;
reg
CUARTlII
;
wire
CUARTOII
;
reg
[
7
:
0
]
CUARTO1I
;
reg
[
1
:
0
]
CUARTOI0
;
reg
[
3
:
0
]
CUARTl11I
;
reg
CUARTOOOl
;
reg
[
8
:
0
]
CUARTIOOl
;
reg
CUARTlOOl
;
reg
[
3
:
0
]
CUARTOIOl
;
reg
CUARTIIOl
;
reg
[
2
:
0
]
CUARTlIOl
;
reg
CUARTOlOl
;
reg
CUARTIlOl
;
reg
CUARTlll
;
reg
CUARTl0l
;
wire
[
1
:
0
]
CUARTllOl
;
wire
[
1
:
0
]
CUARTO0Ol
;
wire
[
3
:
0
]
CUARTI0Ol
;
parameter
CUARTl0Ol
=
0
;
parameter
CUARTO1Ol
=
1
;
parameter
CUARTI1Ol
=
2
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTl1Ol
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTlIOl
<=
3
'b
000
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
CUARTlIOl
[
1
:
0
]
<=
CUARTlIOl
[
2
:
1
]
;
CUARTlIOl
[
2
]
<=
CUARTOl1
;
end
end
end
always
@
(
CUARTlIOl
)
begin
case
(
CUARTlIOl
)
3
'b
000
:
begin
CUARTOOOl
<=
1
'b
0
;
end
3
'b
001
:
begin
CUARTOOOl
<=
1
'b
0
;
end
3
'b
010
:
begin
CUARTOOOl
<=
1
'b
0
;
end
3
'b
011
:
begin
CUARTOOOl
<=
1
'b
1
;
end
3
'b
100
:
begin
CUARTOOOl
<=
1
'b
0
;
end
3
'b
101
:
begin
CUARTOOOl
<=
1
'b
1
;
end
3
'b
110
:
begin
CUARTOOOl
<=
1
'b
1
;
end
default
:
begin
CUARTOOOl
<=
1
'b
1
;
end
endcase
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOOIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTl11I
<=
4
'b
0000
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTOI0
==
CUARTl0Ol
&
(
CUARTOOOl
==
1
'b
1
|
CUARTl11I
==
4
'b
1000
)
)
begin
CUARTl11I
<=
4
'b
0000
;
end
else
begin
CUARTl11I
<=
CUARTl11I
+
1
'b
1
;
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTIOIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTIl1
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTOlOl
==
1
'b
1
)
begin
CUARTIl1
<=
1
'b
1
;
end
end
if
(
CUARTI0I
==
1
'b
1
)
begin
CUARTIl1
<=
1
'b
0
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTlOIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTlI1
<=
1
'b
0
;
end
else
if
(
CUARTIll
==
1
'b
1
)
begin
CUARTlI1
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTIlOl
==
1
'b
1
)
begin
CUARTlI1
<=
1
'b
1
;
end
end
else
begin
CUARTlI1
<=
CUARTlI1
;
end
end
end
assign
CUARTI0Ol
=
CUARTl10
==
1
'b
0
&
CUARTOO1
==
1
'b
0
?
4
'b
0111
:
CUARTl10
==
1
'b
0
&
CUARTOO1
==
1
'b
1
?
4
'b
1000
:
CUARTl10
==
1
'b
1
&
CUARTOO1
==
1
'b
0
?
4
'b
1000
:
4
'b
1001
;
assign
CUARTOl0
=
(
CUARTOI0
==
CUARTl0Ol
)
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOIIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTOI0
<=
CUARTl0Ol
;
CUARTO1I
<=
8
'b
00000000
;
CUARTOlOl
<=
1
'b
0
;
CUARTIlOl
<=
1
'b
0
;
CUARTlI0
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
CUARTOlOl
<=
1
'b
0
;
CUARTlI0
<=
1
'b
0
;
CUARTIlOl
<=
1
'b
0
;
case
(
CUARTOI0
)
CUARTl0Ol
:
begin
if
(
CUARTl11I
==
4
'b
1000
)
begin
CUARTOI0
<=
CUARTO1Ol
;
end
else
begin
CUARTOI0
<=
CUARTl0Ol
;
end
end
CUARTO1Ol
:
begin
if
(
CUARTOIOl
==
CUARTI0Ol
)
begin
CUARTOI0
<=
CUARTI1Ol
;
CUARTOlOl
<=
CUARTIIOl
;
if
(
CUARTIIOl
==
1
'b
0
)
begin
CUARTO1I
<=
{
(
CUARTl10
&
CUARTIOOl
[
7
]
)
,
CUARTIOOl
[
6
:
0
]
}
;
end
end
else
begin
CUARTOI0
<=
CUARTO1Ol
;
end
end
CUARTI1Ol
:
begin
if
(
CUARTl11I
==
4
'b
1110
)
begin
if
(
CUARTOOOl
==
1
'b
0
)
begin
CUARTIlOl
<=
1
'b
1
;
end
end
else
if
(
CUARTl11I
==
4
'b
1111
)
begin
CUARTlI0
<=
1
'b
1
;
CUARTOI0
<=
CUARTl0Ol
;
end
else
begin
CUARTOI0
<=
CUARTI1Ol
;
end
end
default
:
begin
CUARTOI0
<=
CUARTl0Ol
;
end
endcase
end
end
end
assign
CUARTllOl
=
{
CUARTl10
,
CUARTOO1
}
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTIIIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTIOOl
[
8
:
0
]
<=
9
'b
000000000
;
CUARTOIOl
<=
4
'b
0000
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTOI0
==
CUARTl0Ol
)
begin
CUARTIOOl
[
8
:
0
]
<=
9
'b
000000000
;
CUARTOIOl
<=
4
'b
0000
;
end
else
if
(
CUARTl11I
==
4
'b
1111
)
begin
CUARTOIOl
<=
CUARTOIOl
+
1
'b
1
;
case
(
CUARTllOl
)
2
'b
00
:
begin
CUARTIOOl
[
5
:
0
]
<=
CUARTIOOl
[
6
:
1
]
;
CUARTIOOl
[
6
]
<=
CUARTOOOl
;
end
2
'b
11
:
begin
CUARTIOOl
[
7
:
0
]
<=
CUARTIOOl
[
8
:
1
]
;
CUARTIOOl
[
8
]
<=
CUARTOOOl
;
end
default
:
begin
CUARTIOOl
[
6
:
0
]
<=
CUARTIOOl
[
7
:
1
]
;
CUARTIOOl
[
7
]
<=
CUARTOOOl
;
end
endcase
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTlIIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTlOOl
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTl11I
==
4
'b
1111
&
CUARTOO1
==
1
'b
1
)
begin
CUARTlOOl
<=
CUARTlOOl
^
CUARTOOOl
;
end
if
(
CUARTOI0
==
CUARTI1Ol
)
begin
CUARTlOOl
<=
1
'b
0
;
end
end
end
end
assign
CUARTO0Ol
=
{
CUARTl10
,
CUARTIO1
}
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOlIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTll1
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
&
CUARTOO1
==
1
'b
1
&
CUARTl11I
==
4
'b
1111
)
begin
case
(
CUARTO0Ol
)
2
'b
00
:
begin
if
(
CUARTOIOl
==
4
'b
0111
)
begin
CUARTll1
<=
CUARTlOOl
^
CUARTOOOl
;
end
end
2
'b
01
:
begin
if
(
CUARTOIOl
==
4
'b
0111
)
begin
CUARTll1
<=
~
(
CUARTlOOl
^
CUARTOOOl
)
;
end
end
2
'b
10
:
begin
if
(
CUARTOIOl
==
4
'b
1000
)
begin
CUARTll1
<=
CUARTlOOl
^
CUARTOOOl
;
end
end
2
'b
11
:
begin
if
(
CUARTOIOl
==
4
'b
1000
)
begin
CUARTll1
<=
~
(
CUARTlOOl
^
CUARTOOOl
)
;
end
end
default
:
begin
CUARTll1
<=
1
'b
0
;
end
endcase
end
if
(
CUARTOll
==
1
'b
1
)
begin
CUARTll1
<=
1
'b
0
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTIlIl
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTIIOl
<=
1
'b
0
;
CUARTlII
<=
1
'b
1
;
CUARTlll
<=
1
'b
0
;
CUARTl0l
<=
1
'b
0
;
end
else
begin
CUARTlII
<=
1
'b
1
;
CUARTlll
<=
1
'b
0
;
CUARTl0l
<=
1
'b
0
;
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTl10
==
1
'b
1
)
begin
if
(
CUARTOO1
==
1
'b
1
)
begin
if
(
CUARTOIOl
==
4
'b
1001
&
CUARTOI0
==
CUARTO1Ol
)
begin
CUARTlII
<=
1
'b
0
;
CUARTlll
<=
1
'b
1
;
CUARTl0l
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTIIOl
<=
1
'b
1
;
end
end
end
else
begin
if
(
CUARTOIOl
==
4
'b
1000
&
CUARTOI0
==
CUARTO1Ol
)
begin
CUARTlII
<=
1
'b
0
;
CUARTlll
<=
1
'b
1
;
CUARTl0l
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTIIOl
<=
1
'b
1
;
end
end
end
end
else
begin
if
(
CUARTOO1
==
1
'b
1
)
begin
if
(
CUARTOIOl
==
4
'b
1000
&
CUARTOI0
==
CUARTO1Ol
)
begin
CUARTlII
<=
1
'b
0
;
CUARTlll
<=
1
'b
1
;
CUARTl0l
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTIIOl
<=
1
'b
1
;
end
end
end
else
begin
if
(
CUARTOIOl
==
4
'b
0111
&
CUARTOI0
==
CUARTO1Ol
)
begin
CUARTlII
<=
1
'b
0
;
CUARTlll
<=
1
'b
1
;
CUARTl0l
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTIIOl
<=
1
'b
1
;
end
end
end
end
end
if
(
CUARTI0I
==
1
'b
1
)
begin
CUARTIIOl
<=
1
'b
0
;
end
end
end
assign
CUARTOII
=
CUARTIIOl
;
endmodule
