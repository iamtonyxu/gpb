///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: Jabil circuit, Inc.
//
// File: CAN_IF.v
//
// Description: 
//
// CAN Interface Controller
//
// This module provides a CAN (Controller Area Network) interface wrapper for the OPB bus.
// It handles CAN frame transmission and reception for multiple CAN channels, providing
// register-based access to CAN functionality including frame data, control, status,
// and error counting.
//
// Features:
// - 4 CAN channel support (CAN1-4)
// - OPB bus interface for register access
// - Transmit and receive frame handling
// - Error counting and status reporting
//
//
// Targeted device: <Family> <Die> <Package>
// Author: XYL
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

`timescale 1ns / 100ps

module CAN_IF (
    // OPB Interface
    input               OPB_CLK,
    input               OPB_RST,
    input       [31:0]  OPB_DI,
    output      [31:0]  OPB_DO,
    input       [31:0]  OPB_ADDR,

    // GPIO RE/WE Signals
    input               CAN_RE,
    input               CAN_WE,

    // CAN Interface
    output              CAN_TX1,    // CAN BUS, J3, CAN
    output              CAN_TX2,    // CAN BUS, J9, CAND
    output              CAN_TX3,    // CAN BUS, J29/30, CAN_LOC
    output              CAN_TX4,    // CAN BUS, J25, CAN_PEND
    input               CAN_RX1,    // CAN BUS, J3, CAN
    input               CAN_RX2,    // CAN BUS, J9, CAND
    input               CAN_RX3,    // CAN BUS, J29/30, CAN_LOC
    input               CAN_RX4     // CAN BUS, J25, CAN_PEND
);
    // Internal signals for CAN channels
    wire CAN1_RE, CAN1_WE;
    wire CAN2_RE, CAN2_WE;
    wire CAN3_RE, CAN3_WE;
    wire CAN4_RE, CAN4_WE;

    // Output data from CAN channels
    wire [31:0] CAN1_DO;
    wire [31:0] CAN2_DO;
    wire [31:0] CAN3_DO;
    wire [31:0] CAN4_DO;

// Assign RE/WE signals for each CAN channel based on OPB address
    assign CAN1_RE = (OPB_ADDR[14:11] == 4'b0001) && CAN_RE;
    assign CAN1_WE = (OPB_ADDR[14:11] == 4'b0001) && CAN_WE;
    assign CAN2_RE = (OPB_ADDR[14:11] == 4'b0010) && CAN_RE;
    assign CAN2_WE = (OPB_ADDR[14:11] == 4'b0010) && CAN_WE;
    assign CAN3_RE = (OPB_ADDR[14:11] == 4'b0100) && CAN_RE;
    assign CAN3_WE = (OPB_ADDR[14:11] == 4'b0100) && CAN_WE;
    assign CAN4_RE = (OPB_ADDR[14:11] == 4'b1000) && CAN_RE;
    assign CAN4_WE = (OPB_ADDR[14:11] == 4'b1000) && CAN_WE;

// Assign output data from CAN channels to OPB_DO
    assign OPB_DO = (OPB_ADDR[14:11] == 4'b0001) ? CAN1_DO :
                    (OPB_ADDR[14:11] == 4'b0010) ? CAN2_DO :
                    (OPB_ADDR[14:11] == 4'b0100) ? CAN3_DO :
                    (OPB_ADDR[14:11] == 4'b1000) ? CAN4_DO : 32'h00000000;

// CAN1 Interface Instance
CORECAN_wrapper CAN1_inst (
    // OPB Interface
    .OPB_CLK(OPB_CLK),
    .OPB_RST(OPB_RST),
    .OPB_ADDR(OPB_ADDR[10:0]),
    .OPB_DI(OPB_DI),
    .OPB_DO(CAN1_DO),
    .OPB_WE(CAN1_WE),
    .OPB_RE(CAN1_RE),

    // CAN Interface
    .CAN_TX_EN_N(),
    .CAN_TX(CAN_TX1),
    .CAN_RX(CAN_RX1)
);

// CAN2 Interface Instance
CORECAN_wrapper CAN2_inst (
    // OPB Interface
    .OPB_CLK(OPB_CLK),
    .OPB_RST(OPB_RST),
    .OPB_ADDR(OPB_ADDR[10:0]),
    .OPB_DI(OPB_DI),
    .OPB_DO(CAN2_DO),
    .OPB_WE(CAN2_WE),
    .OPB_RE(CAN2_RE),

    // CAN Interface
    .CAN_TX_EN_N(),
    .CAN_TX(CAN_TX2),
    .CAN_RX(CAN_RX2)
);

// CAN3 Interface Instance
CORECAN_wrapper CAN3_inst (
    // OPB Interface
    .OPB_CLK(OPB_CLK),
    .OPB_RST(OPB_RST),
    .OPB_ADDR(OPB_ADDR[10:0]),
    .OPB_DI(OPB_DI),
    .OPB_DO(CAN3_DO),
    .OPB_WE(CAN3_WE),
    .OPB_RE(CAN3_RE),

    // CAN Interface
    .CAN_TX_EN_N(),
    .CAN_TX(CAN_TX3),
    .CAN_RX(CAN_RX3)
);

// CAN4 Interface Instance
CORECAN_wrapper CAN4_inst (
    // OPB Interface
    .OPB_CLK(OPB_CLK),
    .OPB_RST(OPB_RST),
    .OPB_ADDR(OPB_ADDR[10:0]),
    .OPB_DI(OPB_DI),
    .OPB_DO(CAN4_DO),
    .OPB_WE(CAN4_WE),
    .OPB_RE(CAN4_RE),

    // CAN Interface
    .CAN_TX_EN_N(),
    .CAN_TX(CAN_TX4),
    .CAN_RX(CAN_RX4)
);

endmodule

/*
// CoreCan IP generated by Libero
module CORECAN_C0(
    // APB Interface
    input PCLK,
    input PRESETN,
    input PSEL,
    input PENABLE,
    input PWRITE,
    input [10:0] PADDR,
    input [31:0] PWDATA,
    output [31:0] PRDATA,
    output PREADY,
    output INT_N,

    // CAN Interface
    output CAN_TX_EN_N,
    output CAN_TX,
    input CAN_RX
);
*/