//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
`timescale 1ns/100ps
module
UART_UART_0_fifo_256x8
(
CUARTI01
,
CUARTl01
,
CUARTO11
,
CUARTI11
,
WRB
,
RDB
,
RESET
,
FULL
,
EMPTY
)
;
output
[
7
:
0
]
CUARTI01
;
input
CUARTl01
;
input
CUARTO11
;
input
[
7
:
0
]
CUARTI11
;
input
WRB
;
input
RDB
;
input
RESET
;
output
FULL
;
output
EMPTY
;
parameter
[
7
:
0
]
CUARTllII
=
64
;
wire
[
7
:
0
]
CUARTI01
;
wire
FULL
,
EMPTY
;
CUARTO0II
CUARTO0II
(
.CUARTI0OI
(
CUARTI11
)
,
.CUARTl0OI
(
CUARTI01
)
,
.CUARTI0II
(
WRB
)
,
.CUARTl0II
(
RDB
)
,
.CUARTO1II
(
CUARTO11
)
,
.CUARTI1II
(
FULL
)
,
.CUARTl1II
(
EMPTY
)
,
.CUARTOOlI
(
GEQTH
)
,
.CUARTlI
(
RESET
)
,
.CUARTllII
(
CUARTllII
)
)
;
endmodule
module
CUARTO0II
(
CUARTO1II
,
CUARTlI
,
CUARTI0OI
,
CUARTl0II
,
CUARTI0II
,
CUARTllII
,
CUARTl0OI
,
CUARTI1II
,
CUARTl1II
,
CUARTOOlI
)
;
parameter
CUARTIOlI
=
16
;
parameter
CUARTlOlI
=
4
;
parameter
CUARTOIlI
=
8
;
input
CUARTO1II
;
input
CUARTlI
;
input
[
CUARTOIlI
-
1
:
0
]
CUARTI0OI
;
input
CUARTl0II
;
input
CUARTI0II
;
input
[
7
:
0
]
CUARTllII
;
output
[
CUARTOIlI
-
1
:
0
]
CUARTl0OI
;
output
CUARTI1II
;
output
CUARTl1II
;
output
CUARTOOlI
;
wire
CUARTO1II
;
wire
CUARTlI
;
wire
[
CUARTOIlI
-
1
:
0
]
CUARTI0OI
;
wire
CUARTl0II
;
wire
CUARTI0II
;
reg
[
CUARTOIlI
-
1
:
0
]
CUARTl0OI
;
wire
CUARTI1II
;
wire
CUARTl1II
;
wire
CUARTOOlI
;
wire
[
CUARTOIlI
-
1
:
0
]
CUARTIIlI
;
reg
CUARTlIlI
;
reg
[
CUARTlOlI
-
1
:
0
]
CUARTOllI
;
reg
[
CUARTlOlI
-
1
:
0
]
CUARTIllI
;
reg
[
CUARTlOlI
-
1
:
0
]
CUARTlllI
;
assign
CUARTI1II
=
(
CUARTOllI
==
CUARTIOlI
-
1
)
?
1
'b
1
:
1
'b
0
;
assign
CUARTl1II
=
(
CUARTOllI
==
0
)
?
1
'b
1
:
1
'b
0
;
assign
CUARTOOlI
=
(
CUARTOllI
>=
CUARTllII
)
?
1
'b
1
:
1
'b
0
;
always
@
(
posedge
CUARTO1II
or
negedge
CUARTlI
)
begin
if
(
~
CUARTlI
)
begin
CUARTIllI
<=
{
CUARTlOlI
{
1
'b
0
}
}
;
CUARTlllI
<=
{
CUARTlOlI
{
1
'b
0
}
}
;
CUARTOllI
<=
{
CUARTlOlI
{
1
'b
0
}
}
;
end
else
begin
if
(
~
CUARTl0II
)
begin
if
(
CUARTI0II
)
begin
CUARTOllI
<=
CUARTOllI
-
1
;
end
if
(
CUARTIllI
==
CUARTIOlI
-
1
)
CUARTIllI
<=
{
CUARTlOlI
{
1
'b
0
}
}
;
else
CUARTIllI
<=
CUARTIllI
+
1
;
end
if
(
~
CUARTI0II
)
begin
if
(
CUARTOllI
>=
CUARTIOlI
)
begin
$display
(
"\nERROR at time %0t:"
,
$time
)
;
$display
(
"FIFO Overflow\n"
)
;
$stop
;
end
if
(
CUARTl0II
)
begin
CUARTOllI
<=
CUARTOllI
+
1
;
end
if
(
CUARTlllI
==
CUARTIOlI
-
1
)
CUARTlllI
<=
{
CUARTlOlI
{
1
'b
0
}
}
;
else
CUARTlllI
<=
CUARTlllI
+
1
;
end
end
end
always
@
(
posedge
CUARTO1II
or
negedge
CUARTlI
)
begin
if
(
~
CUARTlI
)
begin
CUARTlIlI
<=
1
'b
0
;
end
else
begin
CUARTlIlI
<=
CUARTl0II
;
if
(
CUARTlIlI
==
1
'b
0
)
begin
CUARTl0OI
<=
CUARTIIlI
;
end
else
begin
CUARTl0OI
<=
CUARTl0OI
;
end
end
end
CUARTO0lI
CUARTO0lI
(
.CUARTII
(
CUARTO1II
)
,
.CUARTI0OI
(
CUARTI0OI
)
,
.CUARTl0OI
(
CUARTIIlI
)
,
.CUARTI0lI
(
CUARTlllI
)
,
.CUARTl0lI
(
CUARTIllI
)
,
.CUARTI0II
(
CUARTI0II
)
,
.CUARTl0II
(
CUARTl0II
)
)
;
endmodule
module
CUARTO0lI
(
CUARTII
,
CUARTI0OI
,
CUARTl0lI
,
CUARTI0lI
,
CUARTI0II
,
CUARTl0II
,
CUARTl0OI
)
;
parameter
CUARTO1lI
=
8
;
parameter
CUARTI1lI
=
16
;
parameter
CUARTl1lI
=
4
;
input
CUARTII
;
input
[
CUARTl1lI
-
1
:
0
]
CUARTl0lI
;
input
[
CUARTl1lI
-
1
:
0
]
CUARTI0lI
;
input
CUARTI0II
;
input
CUARTl0II
;
input
[
CUARTO1lI
-
1
:
0
]
CUARTI0OI
;
output
[
CUARTO1lI
-
1
:
0
]
CUARTl0OI
;
wire
[
CUARTl1lI
-
1
:
0
]
CUARTl0lI
;
wire
[
CUARTl1lI
-
1
:
0
]
CUARTI0lI
;
wire
CUARTI0II
;
wire
CUARTl0II
;
reg
[
CUARTO1lI
-
1
:
0
]
CUARTl0OI
;
reg
[
CUARTO1lI
-
1
:
0
]
CUARTOO0I
[
CUARTI1lI
-
1
:
0
]
;
always
@
(
posedge
CUARTII
)
begin
if
(
CUARTI0II
==
1
'b
0
)
begin
CUARTOO0I
[
CUARTI0lI
]
=
CUARTI0OI
;
end
end
always
@
(
posedge
CUARTII
)
begin
if
(
CUARTl0II
==
1
'b
0
)
begin
CUARTl0OI
=
CUARTOO0I
[
CUARTl0lI
]
;
end
end
endmodule
